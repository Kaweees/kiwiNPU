`define FP_WIDTH 16
`define FP_FRACTIONAL 8
